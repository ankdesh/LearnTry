* NMOS Sweep Vds based on image

* Include Sky130 PDK models
.lib "/home/ankdesh/.volare/volare/sky130/versions/0fe599b2afb6708d281543108caf8310912f54af/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* Netlist Description
* Mname drain gate source body model w l
XM1 vdd n1 0 0 sky130_fd_pr__nfet_01v8 w=1 l=0.15
R1 in n1 55
Vdd vdd 0 2.5
Vin in 0 2.5

* Simulation Commands
.control
    dc Vin 0.1 1.8 0.1 Vdd 0 2.5 0.5

    print v(in) i(vdd)
    quit

.endc

.end
