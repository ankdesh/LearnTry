* Sky130 Inverter Simulation

* Include Sky130 PDK models
.lib "/home/ankdesh/.volare/volare/sky130/versions/0fe599b2afb6708d281543108caf8310912f54af/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

.param VDD=1.8

* Power Supply
Vsupply vdd 0 DC VDD

* Input Signal
Vin in 0 PULSE(0 VDD 1ns 100ps 100ps 10ns 20ns)

* Inverter Circuit
* Mname drain gate source body model w l
XM1 out in 0 0 sky130_fd_pr__nfet_01v8 w=1 l=0.15
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 w=2 l=0.15

* Transient Analysis
.tran 0.01ns 40ns

.control
run
plot in out
.endc

.end
