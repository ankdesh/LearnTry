** sch_path: /home/ankdesh/explore/LearnTry/eda/xschem/mos_characterstics/dc_sweep.sch
**.subckt dc_sweep
XM1 vds vgs GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
vgs vgs GND 0
vds vds GND 0
**** begin user architecture code

value=.lib /home/ankdesh/explore/eda/open_pdks/sky130/sky130B/libs.tech/ngspice/sky130.lib.spice tt
.dc vgs 0 1.8 1m vds 0 1.8 0.5
.save all
.end

**** end user architecture code
**.ends
.GLOBAL GND
.end
